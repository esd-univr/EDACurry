.subckt OPAMP1_V1 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1.49918
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V2 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=0.569543
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V3 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=1.018419e-01 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V4 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=2.776686e-05 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V5 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=3.293883e-05 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V6 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=5.511144e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V7 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=5.576174e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V8 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=7.873770e-09 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V9 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=3.200863e-09 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V10 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1.45487
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V11 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=3.682300e-05 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V12 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.295962e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V13 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1.208438e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V14 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=4.485598e-06 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V15 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=3.444165e-09 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V16 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=8.790433e-07 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V17 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=3.758719e-11 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V18 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=4.825449e-06 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V19 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=3.653454e-06 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V20 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=2.912766e-04 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V21 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=0.549312
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V22 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=0.720294
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V23 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=5.976959e-02 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V24 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=1.400570e-11 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V25 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=8.887213e-09 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V26 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=4.682082e-04 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V27 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=1.333397e-11 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V28 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1.09297
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V29 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1.28547
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V30 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=1.378845e-11 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V31 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1.49145
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V32 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=3.574824e-07 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V33 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1.27846
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V34 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=7.288107e-11 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V35 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1.20589
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V36 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.951395e-06 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V37 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1.02678
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V38 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=1.074584e-05 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V39 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=3.686228e-05 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V40 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=9.758466e-11 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V41 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=6.702007e-03 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V42 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=2.322870e-11 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V43 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=1.200885e-11 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V44 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=5.518665e-06 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V45 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=0.96978
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V46 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=0.70694
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V47 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=1.084375e-02 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V48 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=9.871919e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V49 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=1.613495e-02 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V50 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=3.939603e-11 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V51 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=6.129082e-13 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V52 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=8.060952e-07 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V53 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=1.028557e-11 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V54 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=0.524713
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V55 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=1.668147e-05 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V56 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=6.912690e-06 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V57 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=0.582627
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V58 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=2.863590e-05 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V59 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=2.046663e-02 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V60 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=0.878971
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V61 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=7.430938e-07 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V62 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=5.106783e-06 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V63 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=5.344025e-06 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V64 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=1.222466e-05 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V65 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=4.990203e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V66 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=7.243119e-06 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V67 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=8.764756e-02 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V68 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=0.73554
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V69 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=6.076998e-04 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V70 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=4.247870e-07 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V71 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=0.773124
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V72 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=9.825158e-06 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V73 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=5.432734e-06 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V74 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=3.394381e-02 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V75 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=4.927707e-03 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V76 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=8.609820e-02 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V77 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=0.630601
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V78 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=6.352503e-07 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V79 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=3.851245e-02 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V80 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=1.256285e-02 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V81 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=6.456500e-11 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V82 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=2.447550e-11 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V83 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=8.195862e-06 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V84 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=0.8676
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V85 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1.04377
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V86 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=5.832063e-05 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V87 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=7.479026e-05 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V88 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=1.529055e-11 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V89 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=1.725093e-01 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V90 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=9.928185e-13 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V91 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=1.792802e-01 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V92 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=4.672731e-07 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V93 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=0.666556
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V94 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=5.203326e-04 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V95 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=0.622911
.ends

.subckt OPAMP1_V96 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=3.402984e-05 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V97 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=1.516170e-01 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V98 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=3.932320e-05 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V99 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=2.132880e-05 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V100 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=0.657396
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V101 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=9.933075e-13 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V102 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=0.945404
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V103 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=1.014783e-05 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V104 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=1.061011e-11 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V105 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=0.872151
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V106 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=7.837139e-03 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V107 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=1.817329e-05 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V108 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=0.581611
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V109 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=7.613685e-02 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V110 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=0.554538
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V111 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=5.478626e-06 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V112 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=0.851723
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V113 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1.235210e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V114 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=3.791579e-04 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V115 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=3.754661e-06 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V116 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=0.536045
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V117 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1.42012
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V118 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.051319e-06 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V119 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.207740e-06 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V120 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=1.137965e-01 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V121 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1.13904
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V122 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=8.554528e-09 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V123 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=9.608038e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V124 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=7.000588e-06 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V125 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1.16138
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V126 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=5.660475e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V127 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=1.338895e-06 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V128 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=1.824355e-05 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V129 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=1.013227e-01 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V130 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=8.392517e-09 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V131 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=6.761336e-06 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V132 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=9.487543e-05 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V133 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=0.940049
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V134 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.408511e-06 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V135 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=4.913687e-05 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V136 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=0.927815
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V137 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.915395e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V138 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=1.436719e-11 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V139 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.180041e-06 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V140 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=4.715682e-02 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V141 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=2.563291e-11 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V142 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=0.698502
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V143 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=4.205239e-05 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V144 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=4.752184e-11 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V145 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.623603e-06 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V146 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=9.404520e-03 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V147 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=1.285530e-11 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V148 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=2.592381e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V149 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=6.687621e-05 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V150 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=3.750030e-04 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V151 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=7.843264e-07 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V152 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1.12278
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V153 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.709250e-06 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V154 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=2.172073e-06 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V155 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=5.806271e-02 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V156 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=1.258590e-05 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V157 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=1.306635e-11 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V158 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=1.257823e-05 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V159 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=9.373288e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V160 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=5.584796e-09 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V161 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=4.846179e-07 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V162 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=7.814378e-06 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V163 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=6.470619e-09 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V164 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=3.101354e-06 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V165 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=7.450232e-05 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V166 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=0.52174
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V167 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=2.466520e-09 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V168 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=1.273260e-05 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V169 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=5.869310e-06 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V170 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1.08384
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V171 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=0.54716
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V172 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=0.61168
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V173 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=1.048474e-02 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V174 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=4.517647e-06 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V175 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.757018e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V176 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=1.637774e-05 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V177 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=8.291033e-02 M=1
.ends

.subckt OPAMP1_V178 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=5.063104e-07 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V179 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=6.220380e-06 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V180 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=0.958356
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V181 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=0.667479
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V182 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1.49853
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V183 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1.03507
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V184 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=7.558914e-02 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V185 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=7.246966e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V186 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=4.010606e-11 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V187 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=1.214325e-05 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V188 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=6.597214e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V189 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=9.625752e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V190 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.062088e-06 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V191 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=0.837984
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V192 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1.09611
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V193 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=6.030270e-06 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V194 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=6.771246e-02 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V195 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=6.574644e-02 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V196 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=1.150163e-11 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V197 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=8.460242e-02 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V198 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=5.704468e-07 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V199 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=8.122372e-06 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V200 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=7.185948e-02 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V201 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=1.104564e-11 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V202 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=9.085083e-05 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V203 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=6.274464e-02 M=1
.ends

.subckt OPAMP1_V204 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=1.164020e-12 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V205 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1.10273
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V206 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1.430540e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V207 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=1.338754e-05 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V208 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=1.036743e-11 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V209 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=4.007141e-06 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V210 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=1.067635e-05 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V211 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=7.403349e-06 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V212 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=2.327618e-05 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V213 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1.29133
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V214 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=0.983088
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V215 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=8.899218e-13 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V216 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=6.716648e-02 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V217 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4.924310e-06 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V218 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=4.991316e-05 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V219 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=1.759883e-05 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V220 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=3.993171e-05 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V221 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=2.937499e-06 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V222 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=5.924433e-06 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V223 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=2.841027e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V224 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=2.807420e-02 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V225 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1.12986
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V226 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1.47573
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V227 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=9.652668e-02 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V228 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=7.320974e-02 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V229 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1.05438
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V230 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=6.808545e-06 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V231 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=1.376405e-05 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V232 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.979333e-06 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V233 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=1.497153e-05 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V234 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=2.498536e-05 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V235 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=4.355947e-11 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V236 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=8.054062e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V237 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=4.663129e-05 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V238 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=1.802160e-01 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V239 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=1.218686e-05 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V240 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1.40831
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V241 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1.37845
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V242 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=4.724285e-06 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V243 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=5.208866e-06 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V244 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=1.028870e-05 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V245 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=1.210164e-05 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V246 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=8.273753e-06 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V247 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1.11424
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V248 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1.39376
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V249 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=8.935770e-03 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V250 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1.40638
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V251 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=2.400905e-02 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V252 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=9.028149e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V253 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=0.971768
.ends

.subckt OPAMP1_V254 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1.30015
.ends

.subckt OPAMP1_V255 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4.085549e-06 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V256 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=2.510850e-07 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V257 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=5.186034e-04 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V258 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=5.159592e-13 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V259 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=8.597471e-02 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V260 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=6.337165e-07 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V261 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=4.048004e-11 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V262 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1.35263
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V263 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=1.562481e-05 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V264 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=0.879422
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V265 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=1.677291e-02 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V266 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=1.214198e-05 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V267 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=3.474299e-06 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V268 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=6.525909e-06 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V269 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.049225e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V270 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=3.098325e-05 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V271 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=5.427189e-06 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V272 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=7.407890e-06 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V273 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.432896e-06 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V274 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=3.727264e-02 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V275 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=1.142352e-05 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V276 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=1.816559e-02 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V277 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=4.247360e-06 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V278 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.478731e-06 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V279 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=2.991150e-05 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V280 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1.28931
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V281 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=8.050237e-06 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V282 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1.15935
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V283 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=4.405496e-06 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V284 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=1.034596e-05 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V285 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=6.192623e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V286 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=5.101508e-06 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V287 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.450426e-09 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V288 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=7.746517e-06 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V289 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=1.235099e-11 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V290 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1.49606
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V291 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=2.366892e-11 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V292 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=1.778086e-02 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V293 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=9.797350e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V294 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=1.457520e-05 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V295 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=8.035080e-07 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V296 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=3.948983e-11 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V297 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=3.110297e-11 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V298 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1.003441e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V299 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=7.664268e-06 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V300 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=5.376545e-06 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V301 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=8.843880e-06 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V302 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.117434e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V303 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=4.307858e-05 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V304 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=0.688086
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V305 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=1.069627e-04 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V306 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=6.273950e-02 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V307 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.620708e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V308 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=6.765831e-06 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V309 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=1.823849e-11 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V310 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=0.869252
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V311 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=1.088844e-02 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V312 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=5.601257e-06 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V313 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1.25284
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V314 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=1.892340e-05 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V315 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=4.240175e-05 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V316 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.244463e-06 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V317 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=1.316781e-11 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V318 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=5.500725e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V319 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1.34421
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V320 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=0.606732
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V321 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=2.736584e-05 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V322 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=2.090053e-06 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V323 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=4.683843e-13 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V324 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=9.244433e-07 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V325 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=0.973606
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V326 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=4.568853e-07 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V327 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=6.626103e-11 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V328 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=6.462493e-06 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V329 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=0.914763
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V330 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=4.450665e-02 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V331 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=1.323969e-01 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V332 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=0.882944
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V333 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=2.534995e-02 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V334 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1.19911
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V335 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=1.630566e-02 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V336 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=3.484292e-07 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V337 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=7.712731e-06 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V338 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=1.337745e-05 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V339 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=3.255704e-05 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V340 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=4.163396e-11 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V341 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=3.432991e-06 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V342 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=1.697435e-02 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V343 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=4.222933e-07 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V344 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=0.755934
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V345 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=3.749725e-06 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V346 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=0.791167
.ends

.subckt OPAMP1_V347 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=1.162614e-10 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V348 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=5.443045e-07 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V349 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=1.165006e-05 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V350 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.217657e-06 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V351 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=0.74547
.ends

.subckt OPAMP1_V352 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=8.367724e-02 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V353 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=3.635739e-06 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V354 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=4.755810e-07 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V355 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=4.558173e-05 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V356 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=6.007928e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V357 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=1.059467e-05 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V358 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=4.381726e-07 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V359 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=4.306093e-07 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V360 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=5.118067e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V361 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=0.547646
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V362 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.058395e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V363 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=3.550402e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V364 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=3.022953e-06 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V365 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=3.846305e-05 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V366 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1.49707
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V367 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=1.865380e-05 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V368 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=7.586662e-03 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V369 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=4.077332e-13 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V370 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=8.047181e-11 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V371 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=2.584095e-06 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V372 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=2.126845e-02 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V373 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=2.734893e-05 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V374 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=2.610133e-11 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V375 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=5.989049e-07 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V376 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=9.110772e-02 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V377 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=1.471419e-11 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V378 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=0.941652
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V379 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=9.439100e-06 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V380 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=3.620303e-02 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V381 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=5.055239e-03 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V382 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=9.715652e-06 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V383 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=1.766678e-01 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V384 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=1.404388e-02 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V385 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1.41649
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V386 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1.07095
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V387 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=5.972388e-04 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V388 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=0.602164
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V389 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=5.950819e-02 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V390 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=2.881576e-02 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V391 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=1.350742e-01 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V392 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=0.551583
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V393 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=0.514785
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V394 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=5.140214e-04 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V395 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=1.061382e-05 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V396 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=5.164460e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V397 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=9.566353e-06 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V398 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=7.135503e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V399 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=2.348732e-06 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V400 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.133781e-06 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V401 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=4.340562e-05 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V402 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=4.057382e-11 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V403 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=9.685066e-11 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V404 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1.06816
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V405 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=1.505347e-11 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V406 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=1.036987e-11 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V407 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=2.539163e-06 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V408 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.296114e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V409 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=2.099317e-02 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V410 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=9.532255e-06 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V411 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1.45084
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V412 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1.29845
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V413 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=1.352257e-01 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V414 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.877972e-06 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V415 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=3.701037e-05 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V416 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=1.020070e-04 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V417 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=9.805833e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V418 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=7.053982e-11 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V419 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=3.659615e-07 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V420 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=1.179444e-05 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V421 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=1.180656e-10 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V422 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=1.016055e-02 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V423 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=9.815391e-06 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V424 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=4.723307e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V425 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=3.009484e-11 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V426 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=2.575811e-02 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V427 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=1.041110e-12 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V428 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=6.090846e-02 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V429 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=7.378708e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V430 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=1.064152e-12 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V431 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=0.809705
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V432 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=1.280064e-05 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V433 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=1.208252e-05 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V434 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=1.284675e-01 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V435 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=7.677884e-06 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V436 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=4.570455e-05 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V437 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=5.376330e-06 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V438 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=0.601838
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V439 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=1.924939e-06 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V440 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=7.197341e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V441 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=1.453154e-02 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V442 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=1.148508e-05 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V443 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=5.259852e-07 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V444 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=1.227367e-01 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V445 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=0.960213
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V446 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=3.662558e-07 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V447 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=2.753239e-06 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V448 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=1.175787e-12 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V449 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=2.483202e-11 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V450 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.556898e-06 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V451 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=0.874858
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V452 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=1.089556e-02 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V453 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=5.240840e-06 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V454 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.305292e-06 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V455 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=1.114287e-01 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V456 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=9.354487e-06 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V457 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1.100941e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V458 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=5.323563e-06 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V459 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=0.668371
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V460 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=1.203777e-05 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V461 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=1.056254e-05 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V462 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=1.160365e-05 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V463 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=4.299916e-04 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V464 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=4.033043e-03 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V465 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=3.898010e-06 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V466 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=3.761266e-06 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V467 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1.13625
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V468 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=5.741766e-06 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V469 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=3.527781e-05 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V470 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=6.150441e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V471 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=1.498733e-02 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V472 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=3.009689e-11 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V473 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=1.001181e-02 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V474 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1.34393
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V475 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=7.098876e-04 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V476 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=7.233036e-05 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V477 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=1.313614e-10 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V478 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.084647e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V479 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=2.991914e-05 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V480 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1.19853
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V481 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=3.177040e-05 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V482 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=5.400685e-04 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V483 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.889073e-06 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V484 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=0.771674
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V485 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=1.013159e-05 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V486 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1.37182
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V487 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.857485e-06 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V488 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1.44951
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V489 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1.21086
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V490 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=6.583078e-02 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V491 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.817261e-03 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V492 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=0.657702
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V493 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=9.063371e-06 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V494 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=6.521380e-09 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V495 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=9.519078e-06 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V496 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.453906e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V497 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=0.575329
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V498 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=6.441062e-02 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V499 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=2.913855e-11 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V500 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=6.012201e-05 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V501 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=3.662409e-05 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V502 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=4.101405e-05 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V503 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1.0781
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V504 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=1.055484e-02 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V505 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=8.028383e-02 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V506 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=7.913776e-02 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V507 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=4.069049e-09 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V508 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.245683e-06 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V509 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=1.309235e-06 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V510 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=1.743657e-05 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V511 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=7.545367e-09 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V512 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=5.083870e-07 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V513 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=3.506665e-04 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V514 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=7.324414e-06 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V515 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1.2204
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V516 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=0.561906
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V517 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=1.322158e-06 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V518 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1.30873
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V519 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=8.237359e-02 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V520 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=5.490448e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V521 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=4.393660e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V522 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=0.992725
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V523 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=3.992470e-06 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V524 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=7.184333e-06 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V525 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=5.419648e-06 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V526 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=2.100555e-11 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V527 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=2.063426e-01 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V528 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=0.97265
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V529 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=6.717128e-07 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V530 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=2.715369e-06 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V531 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=7.804587e-06 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V532 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=1.442296e-01 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V533 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=8.140382e-02 M=1
.ends

.subckt OPAMP1_V534 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=5.836450e-03 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V535 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=7.224037e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V536 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=1.376563e-05 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V537 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=4.572919e-11 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V538 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=0.735039
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V539 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=1.180877e-01 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V540 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=1.752086e-02 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V541 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=6.820605e-02 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V542 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=5.307392e-11 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V543 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1.382736e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V544 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=0.798099
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V545 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=1.746866e-11 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V546 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=6.034819e-06 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V547 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1.19735
.ends

.subckt OPAMP1_V548 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=9.346357e-05 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V549 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.653522e-06 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V550 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=7.682531e-05 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V551 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=1.101531e-10 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V552 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=5.447745e-09 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V553 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=1.609236e-11 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V554 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=8.959487e-02 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V555 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=5.875288e-07 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V556 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=0.575344
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V557 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=9.419585e-07 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V558 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=0.591934
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V559 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=9.377967e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V560 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=4.235645e-13 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V561 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1.16354
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V562 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=5.705287e-06 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V563 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=1.231355e-05 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V564 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=5.117278e-06 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V565 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1.39352
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V566 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=8.852092e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V567 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.156736e-06 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V568 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=6.021230e-13 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V569 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=3.080734e-09 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V570 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=1.164780e-10 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V571 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=3.382083e-02 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V572 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=4.767862e-06 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V573 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=5.713232e-06 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V574 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1.180657e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V575 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=2.739002e-06 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V576 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=1.180406e-02 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V577 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=6.040284e-06 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V578 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=8.988918e-11 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V579 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1.085886e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V580 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=4.401777e-05 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V581 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=0.651207
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V582 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=9.255719e-06 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V583 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4.736293e-06 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V584 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=4.416906e-07 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V585 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=3.355690e-09 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V586 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=8.746126e-02 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V587 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=1.689318e-05 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V588 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=1.910771e-06 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V589 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=6.383525e-02 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V590 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=1.438290e-02 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V591 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=2.933796e-04 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V592 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=3.140184e-07 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V593 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=2.472164e-06 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V594 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=2.430882e-06 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V595 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=6.622997e-02 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V596 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=6.635975e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V597 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=0.597352
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V598 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=3.327071e-04 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V599 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=3.836026e-06 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V600 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=5.742660e-06 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V601 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1.08237
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V602 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=0.830859
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V603 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1.29854
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V604 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.130137e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V605 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=6.322013e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V606 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=9.538295e-02 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V607 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=5.936623e-02 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V608 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=1.369874e-05 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V609 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=3.723784e-09 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V610 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=9.427185e-06 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V611 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=3.209898e-02 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V612 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=4.194667e-11 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V613 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=9.981837e-06 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V614 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1.3319
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V615 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=5.413431e-06 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V616 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=0.62001
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V617 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=5.852638e-09 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V618 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=0.765066
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V619 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=7.709660e-06 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V620 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=1.666579e-05 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V621 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=1.574590e-05 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V622 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=0.780082
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V623 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=0.735236
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V624 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=5.915917e-06 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V625 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=8.565384e-02 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V626 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.086953e-06 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V627 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=1.547076e-11 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V628 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1.46019
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V629 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=3.293001e-06 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V630 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=1.827782e-11 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V631 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=4.160140e-04 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V632 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=0.514918
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V633 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1.11941
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V634 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=4.353669e-05 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V635 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=3.891782e-06 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V636 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=8.608387e-06 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V637 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=0.78272
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V638 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=5.051325e-02 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V639 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=3.990238e-06 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V640 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=4.063810e-05 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V641 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=6.520845e-05 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V642 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.764985e-06 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V643 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=1.120091e-02 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V644 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=5.641305e-09 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V645 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=9.325422e-07 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V646 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=6.760133e-05 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V647 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=5.891008e-06 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V648 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.067692e-06 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V649 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.990385e-06 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V650 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=7.934993e-11 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V651 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=7.900785e-13 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V652 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=7.272996e-05 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V653 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=1.525966e-05 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V654 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=1.016647e-05 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V655 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=1.470390e-06 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V656 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=3.214018e-06 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V657 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=2.802394e-06 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V658 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=4.512283e-11 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V659 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=4.467068e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V660 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=0.827748
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V661 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=7.269006e-06 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V662 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=5.515418e-06 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V663 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=1.253336e-01 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V664 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=3.085327e-05 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V665 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=4.048660e-06 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V666 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=8.465704e-09 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V667 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=1.158547e-10 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V668 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=3.243043e-05 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V669 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=1.954184e-01 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V670 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=5.215021e-04 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V671 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1.26691
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V672 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=1.476321e-06 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V673 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=4.280929e-02 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V674 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=1.120109e-01 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V675 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=1.354484e-02 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V676 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.526673e-06 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V677 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=2.457693e-02 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V678 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1.39065
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V679 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=7.101631e-04 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V680 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.261957e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V681 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=2.446120e-04 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V682 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=7.915846e-09 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V683 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=2.555577e-07 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V684 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=5.990608e-02 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V685 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1.0409
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V686 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=6.556476e-09 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V687 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=2.078549e-05 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V688 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=3.442609e-06 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V689 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=3.093461e-02 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V690 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=3.466288e-11 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V691 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=3.715928e-09 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V692 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.231563e-06 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V693 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=2.618719e-11 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V694 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=4.004374e-06 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V695 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=2.401218e-11 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V696 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=0.871628
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V697 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=2.825649e-06 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V698 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=6.916409e-06 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V699 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=5.515575e-06 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V700 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=8.377085e-02 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V701 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=0.960932
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V702 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=0.548351
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V703 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=1.105974e-05 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V704 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1.41897
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V705 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1.12768
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V706 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=0.89647
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V707 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=4.672850e-06 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V708 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1.39598
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V709 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=7.482052e-07 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V710 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=2.174020e-07 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V711 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1.26082
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V712 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=3.283198e-06 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V713 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=4.952584e-07 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V714 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=2.154481e-02 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V715 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=5.018921e-05 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V716 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.677701e-09 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V717 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=1.452106e-11 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V718 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=6.412011e-06 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V719 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=1.589884e-02 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V720 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=2.376914e-09 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V721 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=9.304896e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V722 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=0.823604
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V723 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.562389e-06 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V724 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1.25456
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V725 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=9.614434e-06 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V726 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=1.014184e-12 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V727 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=6.371092e-04 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V728 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=6.528067e-02 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V729 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=0.601598
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V730 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=7.274484e-09 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V731 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=1.429618e-11 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V732 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=1.165262e-06 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V733 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=1.390428e-01 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V734 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=6.903588e-13 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V735 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=0.541759
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V736 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=7.582068e-13 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V737 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=5.486189e-02 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V738 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=4.510421e-05 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V739 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1.28594
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V740 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=0.557739
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V741 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=9.749707e-03 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V742 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=1.951224e-06 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V743 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=0.959085
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V744 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=7.554551e-02 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V745 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=4.323174e-06 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V746 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=8.764323e-13 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V747 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=6.429235e-05 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V748 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1.11447
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V749 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=3.687684e-06 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V750 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=6.814085e-09 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V751 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1.11543
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V752 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=5.947719e-06 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V753 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=9.196757e-06 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V754 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=1.953716e-05 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V755 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=0.565811
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V756 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=7.810368e-06 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V757 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=0.856159
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V758 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=8.788768e-07 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V759 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=6.238524e-05 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V760 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=0.873593
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V761 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=5.147005e-06 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V762 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=2.868648e-06 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V763 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=6.364567e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V764 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=3.341638e-06 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V765 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=6.587142e-02 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V766 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=1.400844e-11 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V767 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=1.119057e-11 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V768 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=2.735387e-02 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V769 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=8.252331e-02 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V770 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=4.054600e-11 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V771 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=1.306002e-05 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V772 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=1.153497e-05 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V773 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=2.438454e-02 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V774 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=8.815794e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V775 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=1.171383e-04 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V776 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=4.118174e-07 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V777 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=4.217527e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V778 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=3.669366e-11 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V779 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=8.100796e-03 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V780 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=5.432412e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V781 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=7.073150e-11 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V782 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=4.389253e-04 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V783 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1.17056
.ends

.subckt OPAMP1_V784 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=1.052619e-05 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V785 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=1.040854e-02 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V786 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.595312e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V787 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=2.748348e-11 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V788 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=3.066199e-06 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V789 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.194310e-09 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V790 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=1.513283e-11 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V791 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=4.224580e-04 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V792 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=6.906873e-13 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V793 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=5.873840e-06 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V794 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=0.660514
.ends

.subckt OPAMP1_V795 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1.379182e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V796 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=7.262859e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V797 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=2.850393e-05 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V798 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.394533e-06 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V799 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=4.030548e-02 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V800 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=1.439648e-05 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V801 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=2.926553e-11 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V802 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=6.474781e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V803 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=9.870667e-07 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V804 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=2.020849e-05 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V805 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=4.496220e-06 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V806 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=1.323261e-05 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V807 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=3.477986e-02 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V808 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=2.972508e-06 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V809 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=0.921619
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V810 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=1.840205e-01 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V811 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=5.696321e-04 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V812 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=2.151598e-02 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V813 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=2.162334e-05 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V814 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=4.590654e-07 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V815 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=5.054648e-07 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V816 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.736250e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V817 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=2.474032e-05 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V818 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=0.825819
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V819 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=1.261424e-01 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V820 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=7.677640e-09 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V821 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=2.902410e-05 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V822 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=8.690096e-07 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V823 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=2.449667e-06 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V824 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=5.061783e-02 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V825 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=1.739622e-05 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V826 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=2.077883e-05 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V827 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=1.047884e-02 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V828 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=5.939816e-02 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V829 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=1.684156e-06 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V830 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=9.736165e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V831 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=1.343671e-11 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V832 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=1.142958e-05 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V833 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=8.079714e-06 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V834 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=6.771932e-02 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V835 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=7.539421e-07 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V836 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=6.543944e-06 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V837 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=7.803745e-06 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V838 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=6.156066e-09 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V839 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=3.970012e-06 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V840 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=4.607936e-05 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V841 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=6.512234e-05 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V842 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=2.706008e-05 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V843 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=9.356032e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V844 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=0.744361
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V845 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.337978e-06 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V846 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1.12567
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V847 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=8.523119e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V848 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=1.340682e-05 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V849 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=7.643842e-02 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V850 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=1.410375e-05 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V851 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=8.408120e-02 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V852 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=1.904041e-07 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V853 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1.465448e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V854 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=1.937032e-01 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V855 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=0.893917
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V856 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=0.682669
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V857 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=3.811612e-06 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V858 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=3.181340e-06 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V859 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=7.367995e-06 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V860 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=1.027772e-05 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V861 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=9.422631e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V862 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=0.709989
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V863 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.473556e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V864 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=1.605108e-06 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V865 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=7.059618e-02 M=1
.ends

.subckt OPAMP1_V866 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=5.455796e-11 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V867 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=2.698427e-05 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V868 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=1.004199e-12 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V869 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=0.958361
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V870 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=2.176159e-11 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V871 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=1.380626e-05 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V872 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=8.161452e-02 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V873 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.731630e-06 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V874 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=1.909182e-05 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V875 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=2.216992e-11 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V876 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=6.140974e-02 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V877 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=2.886747e-05 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V878 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=1.960082e-05 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V879 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=8.075829e-03 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V880 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=5.692268e-07 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V881 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=5.819035e-06 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V882 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4.395071e-06 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V883 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=4.322906e-11 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V884 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=1.895793e-05 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V885 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=7.535841e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V886 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=6.660081e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V887 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=1.099689e-05 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V888 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=3.315450e-05 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V889 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=1.176789e-10 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V890 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.074785e-06 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V891 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=0.514249
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V892 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=7.939510e-06 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V893 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=9.559012e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V894 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1.088677e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V895 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1.49596
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V896 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=9.539941e-06 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V897 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=1.340887e-06 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V898 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=1.779680e-05 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V899 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=3.764454e-02 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V900 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=0.921736
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V901 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=4.850418e-07 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V902 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=3.233507e-06 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V903 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=6.962266e-13 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V904 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=0.560235
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V905 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1.15917
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V906 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=4.857194e-11 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V907 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1.19308
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V908 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=2.529243e-06 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V909 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=6.340810e-05 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V910 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=9.542645e-11 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V911 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=0.902488
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V912 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=4.115800e-05 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V913 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=8.640207e-06 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V914 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=1.424802e-11 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V915 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.766171e-06 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V916 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.871379e-06 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V917 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=2.445262e-06 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V918 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=1.112468e-05 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V919 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=7.287391e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V920 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=4.044710e-11 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V921 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=3.089397e-06 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V922 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1.4022
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V923 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=3.244690e-11 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V924 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=8.865269e-02 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V925 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=1.466962e-05 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V926 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=1.549113e-05 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V927 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=7.882826e-06 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V928 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=9.534751e-02 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V929 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=1.479834e-05 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V930 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=6.808643e-02 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V931 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=1.055620e-01 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V932 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=9.126414e-06 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V933 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=4.908102e-06 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V934 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.835204e-09 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V935 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=0.999099
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V936 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=1.086650e-11 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V937 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=2.977328e-05 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V938 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=0.86014
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V939 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=7.483539e-11 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V940 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=2.172017e-11 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V941 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1.36999
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V942 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=9.942908e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V943 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=2.991259e-05 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V944 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=1.021599e-11 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V945 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4.656081e-06 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V946 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=4.970584e-07 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V947 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=4.395093e-05 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V948 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=5.463223e-09 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V949 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=1.207733e-10 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V950 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=3.204775e-06 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V951 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=7.328279e-02 M=1
.ends

.subckt OPAMP1_V952 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=1.187791e-11 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V953 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=1.028800e-05 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V954 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=2.672648e-05 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V955 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=2.826639e-05 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V956 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=6.092282e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V957 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=1.711885e-05 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V958 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=1.063806e-02 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V959 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=5.153374e-07 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V960 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=0.567421
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V961 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1.39462
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V962 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=6.822182e-07 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V963 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=2.129084e-05 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V964 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=6.517289e-09 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V965 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=5.197421e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V966 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=0.505471
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V967 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4.810096e-06 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V968 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=2.971251e-11 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V969 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=1.235211e-05 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V970 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=1.638401e-11 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V971 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=0.921285
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V972 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=1.343527e-01 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V973 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=1.147280e-12 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V974 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=1.287452e-05 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V975 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=9.696408e-03 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V976 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=1.026356e-02 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V977 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=4.298280e-05 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V978 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.619292e-06 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V979 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=9.308894e-02 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V980 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=1.171190e-11 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V981 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=4.759733e-02 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V982 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=4.769437e-05 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V983 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=9.293027e-06 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V984 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=0.522492
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V985 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=1.668971e-05 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V986 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=7.798821e-09 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V987 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=0.770916
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V988 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=0.99085
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V989 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=3.696718e-05 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V990 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=1.410916e-11 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V991 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=1.314264e-05 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V992 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=2.735760e-04 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V993 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.168986e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V994 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=0.795186
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V995 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=5.395193e-11 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V996 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=2.171411e-06 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V997 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=3.075923e-05 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V998 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=1.454756e-05 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V999 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=9.468498e-06 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V1000 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=3.077480e-06 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends
