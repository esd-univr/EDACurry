.subckt OPAMP1_V1 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=9.039958e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V2 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=0.622651
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V3 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=1.134490e-05 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V4 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=4.218444e-06 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V5 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=2.407355e-05 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V6 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1.05249
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V7 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=8.494112e-06 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V8 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=8.218288e-09 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V9 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=6.009316e-09 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V10 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=0.849399
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V11 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=0.556207
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V12 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=0.661904
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V13 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=5.022696e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V14 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1.44069
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V15 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=4.984363e-04 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V16 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=2.711552e-05 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V17 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=8.362018e-02 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V18 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=1.049743e-11 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V19 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=0.551653
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V20 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.285075e-06 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V21 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=8.727410e-13 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V22 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=0.597422
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V23 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.166237e-06 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V24 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=1.582613e-05 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V25 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=7.784762e-02 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V26 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=5.973394e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V27 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=3.040698e-05 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V28 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.847011e-09 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V29 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=8.918330e-02 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V30 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=7.952839e-06 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V31 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=3.589928e-09 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V32 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=2.651711e-05 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V33 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.337570e-06 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V34 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=5.625026e-09 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V35 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=4.049399e-06 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V36 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=9.774651e-03 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V37 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=4.851101e-11 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V38 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=1.585455e-02 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V39 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=1.774535e-02 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V40 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1.150317e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V41 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=4.535304e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V42 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=9.123309e-06 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V43 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=7.140674e-04 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V44 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=0.845645
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V45 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=8.459713e-02 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V46 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=3.400315e-06 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V47 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=1.647490e-11 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V48 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=3.265214e-06 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V49 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=1.002147e-11 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V50 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.824769e-06 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V51 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=0.835806
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V52 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=1.254688e-01 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V53 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=0.951487
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V54 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=3.912395e-02 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V55 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.656268e-09 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V56 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=7.780718e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V57 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=6.779578e-02 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V58 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=1.087056e-12 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V59 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=9.172815e-02 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V60 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=0.688051
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V61 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1.22841
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V62 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=7.574758e-02 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V63 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=4.690081e-02 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V64 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=0.962168
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V65 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=7.493229e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V66 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=8.030438e-06 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V67 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=1.519661e-11 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V68 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=2.013038e-02 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V69 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=1.517619e-05 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V70 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1.07534
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V71 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=6.946649e-11 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V72 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=1.499132e-05 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V73 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=3.885909e-11 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V74 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=3.232102e-02 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V75 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=7.274326e-11 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V76 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=1.423299e-05 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V77 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=5.654071e-05 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V78 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=6.866930e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V79 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1.3659
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V80 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=6.833746e-02 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V81 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=4.036052e-05 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V82 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=0.70448
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V83 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=8.399585e-13 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V84 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=1.009668e-10 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V85 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.903758e-06 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V86 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=3.917922e-11 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V87 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1.32491
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V88 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=0.85011
.ends

.subckt OPAMP1_V89 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=1.312029e-01 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V90 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=6.011104e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V91 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1.14654
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V92 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=1.061917e-11 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V93 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=1.128956e-11 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V94 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=1.212583e-01 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V95 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=2.268703e-05 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V96 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=1.037237e-04 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V97 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=1.099314e-05 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V98 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=4.888743e-11 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V99 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=6.565052e-09 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends

.subckt OPAMP1_V100 inn inp out pd xpd vdda vssa 
xd1 vssa vdda primitive_nwd AREA=6.13907e-9 PJ=476.6e-6 M=1
xi0 vssa net69 primitive_nd AREA=1e-12 PJ=4e-6 M=1
xi3 net51 vdda primitive_pd AREA=790e-15 PJ=3.3e-6 M=1
xr0 vssa vdda net51 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xr1 vdda vdda net69 primitive_rdiffp L=2.1e-6 W=700e-9 M=1
xcc01 net12 out primitive_cpoly AREA=4.7e-9 PERI=453.7e-6 M=1
mnm12 net13 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnm11 net56 net56 vssa vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnb02 net27 net27 net21 vssa nmos1 L=4.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
mnpd1 net21 xpd vssa vssa nmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mn001 out net13 vssa vssa nmos1 L=6.05e-6 W=50e-6 AD=55e-12 AS=55e-12 PD=52.2e-6 PS=52.2e-6 NRD=12e-3 NRS=12e-3 M=1
mnpd2 net13 pd vssa vssa nmos1 L=350e-9 W=5.810533e-06 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mnc01 net13 net69 net12 vssa nmos1 L=7.05e-6 W=4e-6 AD=4.4e-12 AS=4.4e-12 PD=6.2e-6 PS=6.2e-6 NRD=150e-3 NRS=150e-3 M=1
mpb02 net27 net51 net158 vdda pmos1 L=22.05e-6 W=5e-6 AD=5.5e-12 AS=5.5e-12 PD=7.2e-6 PS=7.2e-6 NRD=120e-3 NRS=120e-3 M=1
mppd1 net158 xpd vdda vdda pmos1 L=350e-9 W=6.4e-6 AD=7.04e-12 AS=7.04e-12 PD=8.6e-6 PS=8.6e-6 NRD=93.75e-3 NRS=93.75e-3 M=1
mps11 net31 net158 vdda vdda pmos1 L=6.05e-6 W=20e-6 AD=22e-12 AS=22e-12 PD=22.2e-6 PS=22.2e-6 NRD=30e-3 NRS=30e-3 M=1
mpd11 net56 inn net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mp001 out net158 vdda vdda pmos1 L=6.05e-6 W=80e-6 AD=88e-12 AS=88e-12 PD=82.2e-6 PS=82.2e-6 NRD=7.5e-3 NRS=7.5e-3 M=1
mpd12 net13 inp net31 net31 pmos1 L=4.05e-6 W=30e-6 AD=33e-12 AS=33e-12 PD=32.2e-6 PS=32.2e-6 NRD=20e-3 NRS=20e-3 M=1
mpb01 net158 net158 vdda vdda pmos1 L=6.05e-6 W=10e-6 AD=11e-12 AS=11e-12 PD=12.2e-6 PS=12.2e-6 NRD=60e-3 NRS=60e-3 M=1
.ends
