* AD8304 macromodel
.subckt AD8304
I1	0	IN	DC	1Ua
C1	IN	0	1.0N
E1	2	0	IN	1	3K
V1	1	0	0.5	NPN
Q1	IN	2	0	1u
I2	0	3		NPN
Q2	3	3	0	316.2u
I3	0	4		3
Q3	4	4	0	NPN
.MODEL NPN
E2	5	0	POLY (2)23100,0,0,0,1
E3	6	0	POLY (2)43700,0,0,0,1
E4	7	0	6       5      100K
V2	8	7	0.8
R1	8	9	100
C2	9	0	163P
R2	9	VLOG 4.9K
R3	VLOG 0	1000K
.ends
